`include "apb_mem.v"
`include "apb_tx.sv"
`include "apb_intrf.sv"
`include "apb_gen.sv"
`include "apb_drv.sv"
`include "apb_mon.sv"
`include "apb_scb.sv"
`include "apb_env.sv"
`include "top.sv"
